package avalon_st_tb_pkg;

  `include "generator.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "coverage.sv"

endpackage
